magic
tech scmos
timestamp 1668428488
<< nwell >>
rect -74 54 159 64
rect -74 52 160 54
rect -73 -35 160 52
<< ntransistor >>
rect -57 -71 -53 -61
rect -16 -80 -12 -60
rect 49 -80 53 -60
rect 84 -80 88 -60
rect -16 -136 -12 -116
rect 49 -136 53 -116
rect 84 -136 88 -116
<< ptransistor >>
rect -56 -23 -52 25
rect -18 -23 -14 25
rect 45 -21 55 19
rect 83 -23 87 25
rect 117 -22 121 26
<< ndiffusion >>
rect -61 -71 -57 -61
rect -53 -71 -49 -61
rect -21 -80 -16 -60
rect -12 -80 -8 -60
rect 44 -80 49 -60
rect 53 -80 57 -60
rect 79 -80 84 -60
rect 88 -80 92 -60
rect -21 -136 -16 -116
rect -12 -136 -8 -116
rect 44 -136 49 -116
rect 53 -136 57 -116
rect 79 -136 84 -116
rect 88 -136 92 -116
<< pdiffusion >>
rect -59 15 -56 25
rect -66 6 -56 15
rect -59 -4 -56 6
rect -66 -13 -56 -4
rect -59 -23 -56 -13
rect -52 15 -49 25
rect -52 6 -42 15
rect -52 -4 -49 6
rect -52 -13 -42 -4
rect -52 -23 -49 -13
rect -21 15 -18 25
rect -28 6 -18 15
rect -21 -4 -18 6
rect -28 -13 -18 -4
rect -21 -23 -18 -13
rect -14 15 -8 25
rect -14 6 -2 15
rect -14 -4 -8 6
rect -14 -13 -2 -4
rect -14 -23 -8 -13
rect 42 13 45 19
rect 38 4 45 13
rect 42 -2 45 4
rect 38 -15 45 -2
rect 42 -21 45 -15
rect 55 13 57 19
rect 55 4 63 13
rect 55 -2 57 4
rect 55 -15 63 -2
rect 55 -21 57 -15
rect 80 15 83 25
rect 73 6 83 15
rect 80 -4 83 6
rect 73 -13 83 -4
rect 80 -23 83 -13
rect 87 15 90 25
rect 87 6 97 15
rect 87 -4 90 6
rect 87 -13 97 -4
rect 87 -23 90 -13
rect 114 16 117 26
rect 107 7 117 16
rect 114 -3 117 7
rect 107 -12 117 -3
rect 114 -22 117 -12
rect 121 16 124 26
rect 121 7 131 16
rect 121 -3 124 7
rect 121 -12 131 -3
rect 121 -22 124 -12
<< ndcontact >>
rect -66 -71 -61 -61
rect -49 -71 -42 -61
rect -27 -80 -21 -60
rect -8 -80 -2 -60
rect 38 -80 44 -60
rect 57 -80 63 -60
rect 73 -80 79 -60
rect 92 -80 98 -60
rect -27 -136 -21 -116
rect -8 -136 -2 -116
rect 38 -136 44 -116
rect 57 -136 63 -116
rect 73 -136 79 -116
rect 92 -136 98 -116
<< pdcontact >>
rect -66 15 -59 25
rect -66 -4 -59 6
rect -66 -23 -59 -13
rect -49 15 -42 25
rect -49 -4 -42 6
rect -49 -23 -42 -13
rect -28 15 -21 25
rect -28 -4 -21 6
rect -28 -23 -21 -13
rect -8 15 -2 25
rect -8 -4 -2 6
rect -8 -23 -2 -13
rect 38 13 42 19
rect 38 -2 42 4
rect 38 -21 42 -15
rect 57 13 63 19
rect 57 -2 63 4
rect 57 -21 63 -15
rect 73 15 80 25
rect 73 -4 80 6
rect 73 -23 80 -13
rect 90 15 97 25
rect 90 -4 97 6
rect 90 -23 97 -13
rect 107 16 114 26
rect 107 -3 114 7
rect 107 -22 114 -12
rect 124 16 131 26
rect 124 -3 131 7
rect 124 -22 131 -12
<< psubstratepcontact >>
rect -27 -107 -21 -101
rect -83 -161 -73 -152
rect -65 -161 -55 -152
rect -40 -162 -30 -153
rect -17 -163 -7 -154
rect 39 -161 49 -152
rect 61 -161 71 -152
rect 79 -162 89 -153
rect 99 -162 109 -153
<< nsubstratencontact >>
rect -69 45 -59 54
rect -51 45 -41 54
rect -27 45 -17 54
rect -5 45 5 54
rect 33 46 43 55
rect 55 45 65 54
rect 76 44 86 53
rect 95 45 105 54
rect 119 45 129 54
<< polysilicon >>
rect -56 29 -53 33
rect -56 25 -52 29
rect -18 25 -14 37
rect 83 28 86 33
rect 117 30 120 35
rect 83 25 87 28
rect 117 26 121 30
rect 45 19 55 24
rect -56 -27 -52 -23
rect -18 -27 -14 -23
rect -54 -31 -52 -27
rect -17 -32 -14 -27
rect 45 -25 55 -21
rect 45 -30 54 -25
rect 83 -27 87 -23
rect 117 -26 121 -22
rect 84 -32 87 -27
rect -18 -33 -14 -32
rect -15 -54 -12 -50
rect 51 -54 53 -50
rect 85 -54 88 -50
rect -57 -61 -53 -56
rect -16 -60 -12 -54
rect 49 -60 53 -54
rect 84 -60 88 -54
rect -57 -75 -53 -71
rect -57 -79 -54 -75
rect -16 -85 -12 -80
rect 49 -85 53 -80
rect -16 -89 -13 -85
rect 49 -89 52 -85
rect 84 -89 88 -80
rect -16 -116 -12 -110
rect 50 -113 53 -109
rect 85 -113 88 -109
rect 49 -116 53 -113
rect 84 -116 88 -113
rect -16 -139 -12 -136
rect 49 -139 53 -136
rect -16 -143 -13 -139
rect 49 -143 52 -139
rect 84 -142 88 -136
rect -16 -147 -12 -143
rect -16 -151 -13 -147
rect -16 -152 -12 -151
<< polycontact >>
rect -53 29 -49 33
rect 86 28 91 33
rect 120 30 127 35
rect -59 -31 -54 -27
rect -22 -32 -17 -27
rect 54 -30 59 -25
rect 79 -32 84 -27
rect -19 -54 -15 -50
rect 46 -54 51 -50
rect 80 -54 85 -50
rect -54 -79 -50 -75
rect -13 -89 -8 -85
rect 52 -89 57 -85
rect 46 -113 50 -109
rect 81 -113 85 -109
rect -13 -143 -8 -139
rect 52 -143 57 -139
rect -13 -151 -8 -147
<< metal1 >>
rect -73 54 33 55
rect -73 45 -69 54
rect -59 45 -51 54
rect -41 45 -27 54
rect -17 45 -5 54
rect 5 46 33 54
rect 43 54 160 55
rect 43 46 55 54
rect 5 45 55 46
rect 65 53 95 54
rect 65 45 76 53
rect -73 44 76 45
rect 86 45 95 53
rect 105 45 119 54
rect 129 45 160 54
rect 86 44 160 45
rect -73 43 160 44
rect -66 25 -59 43
rect -49 29 -32 33
rect -64 -31 -59 -27
rect -49 -61 -42 -23
rect -37 -27 -32 29
rect -28 25 -21 43
rect 38 19 42 43
rect 73 36 104 40
rect 73 25 80 36
rect 91 28 95 33
rect -37 -32 -22 -27
rect -37 -54 -19 -50
rect -66 -151 -61 -71
rect -37 -75 -33 -54
rect -8 -60 -2 -23
rect 57 -25 63 -21
rect 59 -27 63 -25
rect 59 -30 79 -27
rect 57 -32 79 -30
rect 100 -28 104 36
rect 107 26 114 43
rect 127 30 134 35
rect 124 -28 131 -22
rect 100 -32 131 -28
rect -50 -79 -33 -75
rect 30 -54 46 -50
rect -27 -101 -21 -80
rect 30 -85 34 -54
rect 57 -60 63 -32
rect -8 -89 34 -85
rect 66 -54 80 -50
rect -21 -107 -2 -101
rect 38 -102 44 -80
rect 66 -85 70 -54
rect 57 -89 70 -85
rect 73 -94 79 -80
rect 73 -99 98 -94
rect 38 -106 63 -102
rect -8 -116 -2 -107
rect 18 -113 46 -109
rect -27 -151 -21 -136
rect 18 -139 22 -113
rect 57 -116 63 -106
rect -8 -143 22 -139
rect 66 -113 81 -109
rect 38 -151 44 -136
rect 66 -139 70 -113
rect 92 -116 98 -99
rect 57 -143 70 -139
rect 73 -151 79 -136
rect -86 -152 -21 -151
rect -86 -161 -83 -152
rect -73 -161 -65 -152
rect -55 -153 -21 -152
rect -55 -161 -40 -153
rect -86 -162 -40 -161
rect -30 -154 -21 -153
rect 38 -152 147 -151
rect 38 -154 39 -152
rect -30 -162 -17 -154
rect -86 -163 -17 -162
rect -7 -161 39 -154
rect 49 -161 61 -152
rect 71 -153 147 -152
rect 71 -161 79 -153
rect -7 -162 79 -161
rect 89 -162 99 -153
rect 109 -162 147 -153
rect -7 -163 147 -162
<< metal2 >>
rect -2 -53 16 -44
rect 7 -147 16 -53
rect -13 -151 16 -147
<< labels >>
rlabel metal1 20 47 20 47 1 Vdd
rlabel metal1 16 -158 16 -158 1 gnd
rlabel metal1 -37 29 -37 33 1 Vbiasb
rlabel metal1 14 -89 14 -85 1 Vbias3
rlabel metal1 134 30 134 35 1 Vbias1
rlabel metal1 95 28 95 33 1 Vbias2
<< end >>
